/* tb_lab7_g41_p3.sv
* Hazırlayanlar: Berat Kızılarmut, Ömer Emre Polat
* Notlar: Modül birleştirme testbench */
`timescale 1ns/1ps
module tb_lab7_g41_p3();
logic clk, reset;
logic [31:0] komut;
logic [6:0] opcode;
logic [3:0] aluop;
logic [31:0] rs1_data;
logic [31:0] rs2_data;
logic [31:0] imm;
logic hata;
logic we;
logic [31:0] rd_data;

lab7_g41_p3 dut0(.clk(clk), .reset(reset), .komut(komut), .opcode(opcode), .aluop(aluop), .rs1_data(rs1_data), .rs2_data(rs2_data), .imm(imm), .hata(hata), .we(we), .rd_data(rd_data));
always
begin
    clk = 1; #5;
    clk = 0; #5;
end
initial 
begin
    we = 1; reset = 0;
    rd_data = 32'd1; #10;
    komut = 32'b0100000_10100_00110_001_10011_0000001; #10;
    rd_data = 32'd2; #10;
    komut = 32'b0100000_10100_00110_001_10011_0000001; #10;
    rd_data = 32'd3; #10;
    komut = 32'b010000010100_00110_001_10011_0000011; #10;
    rd_data = 32'd4; #10;
    komut = 32'b000000001011_11001_001_10111_0000011; #10;
    rd_data = 32'd5; #10;
    komut = 32'b01000001010000110001_10011_0000111; #10;
    rd_data = 32'd6; #10;
    komut = 32'b00000000101111001001_10111_0000111; #10;
    rd_data = 32'd7; #10;
    komut = 32'b0100000_10100_00110_001_10011_0001111; #10;
    rd_data = 32'd8; #10;
    komut = 32'b0000000_01011_11001_001_10111_0001111; #10;
    we = 0; reset = 0; rd_data = 32'd1;
    /////////////////R///////////////////////
    komut = 32'b0100000_10100_00110_001_10011_0000001; #10;
    komut = 32'b0100000_10100_00110_001_10011_0000001; #10;
    komut = 32'b0000000_10010_10001_101_11111_0000001; #10;
    komut = 32'b0100000_01110_10101_100_01100_0000001; #10;
    /////////////////I///////////////////////
    komut = 32'b010000010100_00110_001_10011_0000011; #10;
    komut = 32'b000000001011_11001_001_10111_0000011; #10;
    komut = 32'b000000010010_10001_101_11111_0000011; #10;
    komut = 32'b010000001110_10101_100_01100_0000011; #10;
    /////////////////U///////////////////////
    komut = 32'b01000001010000110001_10011_0000111; #10;
    komut = 32'b00000000101111001001_10111_0000111; #10;
    komut = 32'b00000001001010001101_11111_0000111; #10;
    komut = 32'b01000000111010101100_01100_0000111; #10;
    /////////////////B///////////////////////
    komut = 32'b0100000_10100_00110_001_10011_0001111; #10;
    komut = 32'b0000000_01011_11001_001_10111_0001111; #10;
    komut = 32'b0000000_10010_10001_101_11111_0001111; #10;
    komut = 32'b0100000_01110_10101_100_01100_0001111; #10;
    /////////////////HATA////////////////////
    komut = 32'b0100000_10100_00110_001_10011_0010001; #10;
    komut = 32'b0000000_01011_11001_001_10111_0100001; #10;
    komut = 32'b0000000_10010_10001_101_11111_0001001; #10;
    komut = 32'b0100000_01110_10101_100_01100_0101101; #10;
    $stop;
end
endmodule
